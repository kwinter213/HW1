//Hw1, 9/15/17, Originally written by Ben Hill

// Simple Verilog test
module hello_test ();
initial begin
    $display("Hello, CompArch!");
end
endmodule